component traffic_light.CDiagMessage

endpoints {
    dmessage : traffic_light.IDiagMessage
}