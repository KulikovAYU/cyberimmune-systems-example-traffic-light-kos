component traffic_light.CControlSystem

endpoints {
    mode : traffic_light.ControlSystem
}